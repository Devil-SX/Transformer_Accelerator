`include "Types.sv"

module Skew(
    input clk,
    input rst_n,

    input `SINGLE data_in[`SYS_ARRAY_LEN],
    input logic data_valid,
    output Scalar scalar_out[`SYS_ARRAY_LEN], 
);




endmodule