`include "Types.sv"

module #(parameter LENGTH = 1) ShiftedReg(
    input clk,
    input rst_n,
    
);


endmodule