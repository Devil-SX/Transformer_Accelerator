module CIMCore(
    input clk,
    input rst_n,

    
);



endmodule