`ifndef FIXED_SV
`define FIXED_SV

`include "../Types.sv"


`endif